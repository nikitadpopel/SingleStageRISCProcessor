li s1, 0x0004       01101 000 001 00100
sll s1, s1, 4       00111 001 001 00100

li s2, 0x0010       01101 000 010 10000
sll s2, s2, 8       00111 010 010 01000
addi s2, s2, 0x0010 01110 010 010 10000

li s3, 0x000F       01101 000 011 01111

li s4, 0x000F       01101 000 100 01111
sll s4, s4, 4       00111 100 100 00100

li s6, 0x0010       01101 000 110 10000

li s7, 0x0005       01101 000 111 00101


li s0, 0x0001       01101 000 000 00001
sll s0, s0, 8       00111 000 000 01000
addi s0, s0, 0x0001 01110 000 000 00001
sw s0, s6           01011 110 000 00000

addi s0, s0, 0x000F 01110 000 000 01111
sw s0, s6 0x0002    01011 110 000 00010

srl s0, s0, 4       01000 000 000 00100
sw s0, s6, 0x0004   01011 110 000 00100

li s0, 0x000F       01101 000 000 01111
sll s0, s0, 4       00111 000 000 00100
sw s0, s6, 0x0006   01011 110 000 00110

addi s0, s0, 0x000F 01110 000 000 01111
sw s0, s6, 0x0008   01011 110 000 01000
